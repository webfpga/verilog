module fpga_top;
    // instantiate one of these modules:

    // control fade(/*...*/);
    // control rainbow(/*...*/);
    control simple(/*...*/);
    // control random(/*...*/);
endmodule
