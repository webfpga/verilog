//////////////////////////////////////////////////////////////////////
//   ROM holding rainbow colors.  ROM will be made out of a BRAM.
//
module WF_neo_fading_rom ( rd_data, rd_addr,clk);
  output [15:0]  rd_data;
  input   [7:0]  rd_addr;
  input          clk;

  wire [15:0] rd_data1;
  wire [15:0] rd_data;

  // bit reverse ROM data for LSB being brightest.
  assign rd_data = {rd_data1[15],
                    rd_data1[10],rd_data1[11],rd_data1[12],rd_data1[13],rd_data1[14],
                    rd_data1[5],rd_data1[6],rd_data1[7],rd_data1[8],rd_data1[9],
                    rd_data1[0],rd_data1[1],rd_data1[2],rd_data1[3],rd_data1[4]};

                 SB_RAM256x16  ram ( .WDATA(16'b0),
                               .MASK(16'b0),
                               .WADDR(8'b0),
                               .WE(1'b0),
                               .WCLKE(1'b0),
                               .WCLK(1'b0),
                               .RDATA(rd_data1),
                               .RADDR(rd_addr),
                               .RE(1'b1),
                               .RCLKE(1'b1),
                               .RCLK(clk));

defparam ram.INIT_0 = 256'b0001011101000000000101110100000000010011010000000001001101100000000100110110000000001111011000000000111110000000000011111000000000001011101000000000101110100000000001111010000000000111110000000000011111000000000000111100000000000011111000000000001111100000;
defparam ram.INIT_1 = 256'b0010111010000000001011101000000000101010100000000010101010100000001010101010000000100110101000000010011011000000001001101100000000100010111000000010001011100000000111101110000000011111000000000001111100000000000110110000000000011011001000000001101100100000;
defparam ram.INIT_2 = 256'b0100010111000000010001011100000001000001110000000100000111100000010000011110000000111101111000000011111000000000001111100000000000111010001000000011101000100000001101100010000000110110010000000011011001000000001100100100000000110010011000000011001001100000;
defparam ram.INIT_3 = 256'b0101110100000000010111010000000001011001000000000101100100100000010110010010000001010101001000000101010101000000010101010100000001010001011000000101000101100000010011010110000001001101100000000100110110000000010010011000000001001001101000000100100110100000;
defparam ram.INIT_4 = 256'b0111010001000000011101000100000001110000010000000111000001100000011100000110000001101100011000000110110010000000011011001000000001101000101000000110100010100000011001001010000001100100110000000110010011000000011000001100000001100000111000000110000011100000;
defparam ram.INIT_5 = 256'b0110110000000011011100000000001101110000000000110111010000000010011101000000001001110100000000010111100000000001011110000000000101111000000000000111110000000000011111000000000001111100000000000111110000000000011110000000000001111000001000000111100000100000;
defparam ram.INIT_6 = 256'b0101010000001001010110000000100101011000000010010101110000001000010111000000100001011100000001110110000000000111011000000000011101100000000001100110010000000110011001000000011001101000000001010110100000000101011010000000010001101100000001000110110000000100;
defparam ram.INIT_7 = 256'b0011110000001111010000000000111101000000000011110100010000001110010001000000111001000100000011010100100000001101010010000000110101001000000011000100110000001100010011000000110001010000000010110101000000001011010100000000101001010100000010100101010000001010;
defparam ram.INIT_8 = 256'b0010010000010101001010000001010100101000000101010010110000010100001011000001010000101100000100110011000000010011001100000001001100110000000100100011010000010010001101000001001000111000000100010011100000010001001110000001000000111100000100000011110000010000;
defparam ram.INIT_9 = 256'b0000110000011011000100000001101100010000000110110001010000011010000101000001101000010100000110010001100000011001000110000001100100011000000110000001110000011000000111000001100000100000000101110010000000010111001000000001011000100100000101100010010000010110;
defparam ram.INIT_A = 256'b0000000000111101000000000011111000000000001111100000000000011110000000000001111100000000000111110000000000011111000000000001111100000000000111100000010000011110000001000001111000001000000111010000100000011101000010000001110000001100000111000000110000011100;
defparam ram.INIT_B = 256'b0000000011110111000000001111100000000000111110000000000011011000000000001101100100000000110110010000000010111010000000001011101000000000100110100000000010011011000000001001101100000000011110110000000001111100000000000111110000000000010111010000000001011101;
defparam ram.INIT_C = 256'b0000000110110001000000011011001000000001101100100000000110010010000000011001001100000001100100110000000101110100000000010111010000000001010101000000000101010101000000010101010100000001001101010000000100110110000000010011011000000001000101110000000100010111;
defparam ram.INIT_D = 256'b0000001001101011000000100110110000000010011011000000001001001100000000100100110100000010010011010000001000101110000000100010111000000010000011100000001000001111000000100000111100000001111011110000000111110000000000011111000000000001110100010000000111010001;
defparam ram.INIT_E = 256'b0000001100100101000000110010011000000011001001100000001100000110000000110000011100000011000001110000001011101000000000101110100000000010110010000000001011001001000000101100100100000010101010010000001010101010000000101010101000000010100010110000001010001011;
defparam ram.INIT_F = 256'b0000001111100000000000111110000000000011111000000000001111000000000000111100000100000011110000010000001110100010000000111010001000000011100000100000001110000011000000111000001100000011011000110000001101100100000000110110010000000011010001010000001101000101;


  endmodule

